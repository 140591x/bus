`timescale 1ns / 1ps

module tb_ahb_master; 
 
wire HBUSREQ,HLOCK,HWRITE; 
wire [1:0]HTRANS,HSEL; 
wire [31:0]HADDR,HWDATA; 
wire [2:0]HSIZE,HBURST; 
 
reg HGRANT,HREADY,HCLK,HRESETn,BUSREQ,ADDREQ,WRITE,htrans_comp; 
reg [1:0]HRESP; 
reg [31:0]HRDATA; 
reg [1:0]TRANS,SEL; 
reg [31:0]ADDR,WDATA; 
reg [2:0]SIZE,BURST; 
 
ahb_master mst(.HBUSREQ(HBUSREQ),.HLOCK(HLOCK),.HTRANS(HTRANS),.HADDR(HADDR),.HWRITE(HWRITE),.HSIZE(HSIZE),.HBURST(HBURST),.HWDATA(HWDATA),.HSEL(HSEL),.HRESETn(HRESETn),.HCLK(HCLK),.HGRANT(HGRANT),.HREADY(HREADY),.HRESP(HRESP),.HRDATA(HRDATA),.BUSREQ(BUSREQ),.ADDREQ(ADDREQ),.WRITE(WRITE),.ADDR(ADDR),.SIZE(SIZE),.BURST(BURST),.SEL(SEL),.TRANS(TRANS),.WDATA(WDATA)); 
//ahb_master(HBUSREQ,HLOCK,HTRANS,HADDR,HWRITE,HSIZE,HBURST,HWDATA,HSEL,hcount,HRESETn,HCLK,HGRANT,HREADY,HRESP,HRDATA,BUSREQ,ADDREQ,WRITE,ADDR,SIZE,BURST,SEL,TRANS,WDATA); 
initial 
begin 
 HRESETn = 1'b0; 
 HGRANT = 1'b0; 
 HREADY = 1'b0; 
 HCLK = 1'b0; 
 BUSREQ = 1'b0; 
 ADDREQ = 1'b0; 
 WRITE = 1'b0; 
 ADDR=32'h00000000; 
 WRITE=1'b0; 
 SIZE=3'b000; 
 BURST=3'b000; 
 SEL=2'b00; 
 TRANS=2'b00; 
 HRESP = 2'b00; 
 htrans_comp = 1'b0; 
end 
 
always  
#5  HCLK = ~HCLK; 
 
initial 
begin 
#20 HRESETn = 1'b1; 
#5 BUSREQ = 1'b1; 
//WRITE TRANSFER 
//NON SEQ 
#10 BUSREQ = 1'b0;HGRANT = 1'b1;ADDREQ=1'b1;ADDR=32'h00abcdef;WRITE=1'b1;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b00;WDATA=32'hf0f0f0f0; 
#10 ADDREQ = 1'b0; 
#10 HREADY = 1'b1;HRESP = 2'b00; 
//SEQUENTIAL 
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'b11111111111111110000000010101100;WRITE=1'b1;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b01;WDATA=32'b00001111000011110000111100001111; 
#10 ADDREQ = 1'b0;WDATA=32'b10101010101010101010101010101010; 
#10 WDATA=32'b11111111111111110000000010101100; 
#10 WDATA=32'b11001100110011001100110011001100; 
#10 WDATA=32'b10101010101010101010101010101010; 
#10 HREADY = 1'b1;HRESP = 2'b01; 
//IDLE 
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'hbcdabcdb;WRITE=1'b1;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b10;WDATA=32'h0f0f0f0f; 
#10 HREADY = 1'b1;ADDREQ = 1'b0;WDATA=32'haaaaaaaa;HRESP = 2'b00; 
//BUSY  
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'b11111111111111110000000010101100;WRITE=1'b1;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b11;WDATA=32'hfa0f000a; 
#10 ADDREQ = 1'b0;WDATA=32'haaaaaaaa; 
#10 WDATA=32'habcdefac; 
#10 WDATA=32'h09acbdba; 
#10 WDATA=32'hbbbbbbbb; 
#10 HREADY = 1'b1;HRESP = 2'b00; 
#10 HREADY = 1'b0;WDATA=32'hffaaffbb; 
#10 WDATA = 32'hababcdcd; 
#10 WDATA = 32'hcdcdabab; 
#10 HREADY = 1'b1;HRESP = 2'b01; 
#10 HREADY = 1'b0;TRANS = 2'b10;  // time = 245 
//READ TRANSFER 
//NON SEQ 
#10 BUSREQ = 1'b0;HGRANT = 1'b1;ADDREQ=1'b1;ADDR=32'h00001111;WRITE=1'b0;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b00;HRESP = 2'b00; 
#10 ADDREQ = 1'b0;HRDATA = 32'h50505050; 
#10 HREADY = 1'b1; 
//SEQUENTIAL 
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'h00000101;WRITE=1'b0;SIZE=3'b010;BURST=3'b000;SEL=2'b10;TRANS=2'b01; 
#10 ADDREQ = 1'b0;HRDATA = 32'h45454545; 
#10 HRDATA=32'h86868686; 
#10 HRDATA=32'h75757575; 
#10 HRDATA=32'h99994444; 
#10 HREADY = 1'b1; 
//IDLE 
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'hbcdabcdb;WRITE=1'b1;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b10; 
#10 HREADY = 1'b1;ADDREQ = 1'b0;HRDATA=32'haaaaaaaa; 
//BUSY  
#10 HREADY = 1'b0;ADDREQ=1'b1;ADDR=32'h00001111;WRITE=1'b0;SIZE=3'b010;BURST=3'b111;SEL=2'b10;TRANS=2'b11; 
#10 ADDREQ = 1'b0;HRDATA=32'haaaaaaaa; 
#10 HRDATA=32'habcdefac; 
#10 HRDATA=32'h09acbdba; 
#10 HRDATA=32'hbbbbbbbb; 
#10 HREADY = 1'b1; 
#10 HREADY = 1'b0;HRDATA=32'hffaaffbb; 
#10 HRDATA = 32'hababcdcd; 
#10 HRDATA = 32'hcdcdabab; 
#10 HREADY = 1'b1; 
#10 HREADY = 1'b0;TRANS = 2'b10;  // time = 245 
#10 HGRANT = 1'b0;htrans_comp = 1'b1; 
end  
 
endmodule 